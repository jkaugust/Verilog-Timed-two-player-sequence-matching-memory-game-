module GameController();
input Clk,Rst;
output
always @(posedge Clk)
if
