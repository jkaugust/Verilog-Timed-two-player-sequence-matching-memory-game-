//Course Number:6370
//Author: Justin K Augustine 2199
module AccessControl(P,V,Allow,Clk,Rst);
 input P,V,Clk,Rst;
 output Allow;
 reg Allow;
 reg Flag;
 reg [2:0]State;
 parameter INIT=0,B1=1,B2=2,B3=3,B4=4,B5=5,VALID=6;
always@(posedge Clk)
 begin
  if(Rst==1)
  begin
   case(State)
    INIT:
     begin
    Allow<=1'b0;
     if(V==1)     
      begin
       Flag<=0;
       if(P!=1)
        begin
         Flag<=1'b1;
        end
       State<=B1;
      end
     else
      begin
       State<=INIT;
      end  
    end
   B1:
    begin
      if(V==1)
       begin
        if(P!=1)
         begin
         Flag<=1'b1;
         end
        State<=B2;
       end
       else
     begin
     State<=B1;
     end
    end
  B2:
   begin
    if(V==1)
     begin
      if(P!=1)
       begin
        Flag<=1'b1;
       end
       State<=B3;
      end
      else
       begin
       State<=B2;
       end
    end
  B3:
   begin
     if(V==1)
      begin
      if(P!=1)
       begin
        Flag<=1'b1;
       end
      State<=B4;
     end
    else
    begin
     State<=B3;
     end
    end
  B4:
   begin
     if(V==1)
      begin
      if(P!=1)
        begin
         Flag<=1'b1;
        end
      State<=B5;
      end
      else
       begin
        State<=B4;
       end
   end   
   B5:
    begin
     if(V==1)
      begin
       if(P!=1)
        begin
        Flag<=1'b1;
        end
       State<=VALID;
      end 
      else
       begin
        State<=B5;
       end
    end
   VALID:
    begin
     if(Flag==0)
      begin
       Allow<=1'b1;
      end
     else
      begin
       Allow<=1'b0; 
      end
      State<=VALID;
    end
   endcase
 end
 else
  if(Rst==0)
   begin
   State<=INIT;
   end
   else
  begin
   Allow<=1'b0;
   Flag<=1'b0;
   end
end
endmodule
